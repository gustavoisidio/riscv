library verilog;
use verilog.vl_types.all;
entity simulacao32 is
end simulacao32;
