library verilog;
use verilog.vl_types.all;
entity UP is
    port(
        clock           : in     vl_logic;
        reset           : in     vl_logic
    );
end UP;
